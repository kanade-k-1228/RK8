///////////////////////////////////////////////////////////////////////////////////////////////////
// Parallel_ROM ///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                               //
// アドレスの変化を検出したら、ROMにアクセスして、データを取り出す。                             //
//                                                                                               //
//               _   _   _   _   _   _   _   _   _   _   _   _   _   _   _   _   _   _   _   _   //
//  clk        :  |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_| |_ //
//                  :                               :                               :   :        //
//  addr       :  0xXXXX | - - - - - - - - - - - - - : - - - - - - - - - - - - - - - : - : - - - //
//                 _:___                            :                               :   :        // 
//  addr_valid : _| :   |___________________________:_______________________________:___:_______ //
//               ___^ pos clk & valid -> send       :                               :   ;_______ //
//  addr_ready :    |_______________________________:_______________________________:___|        //
//                  :                               :                               :   ;        //
//  mode       :    | sending                       | receiving                     |end| waiting//
//                  :                               :                               :   :        //
//  count      :  - | 0 | 1 | 2 | 3 | 4 | : |62 |63 | 0 | 1 | 2 | 3 | 4 | : |62 |63 |   ;        //
//                  :                               :                               :___:        //
//  data_valid : ___:_______________________________:_______________________________|   |_______ //
//                  :                               :                               :   :        //
//  data       :  PREV_DATA - - - - - - - - - - - - : - | - - - | - - - | - - - | 0x0123_4567    //
//                  :    ___     ___     ___     ___:    ___     ___     ___     ___:   :        //
//  SCL        : ___:___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___:_______ //
//                  :                               :                               :   :        //
//  MOSI       :  - | [31]  | [30]  |   :   |  [0]  |                               |   :        //
//                  :                               :                               :   :        //
//  MISO       :    :                               : [31]  | [30]  |   :   |  [0]  |   :        //
//            [R]  [A] [B] [C]                     [D] [E] [F]                     [G] [H]       //
///////////////////////////////////////////////////////////////////////////////////////////////////


module Parallel_ROM (
    input  logic [23:0] addr,
    output logic [31:0] data,
    output logic        valid
);




endmodule
